module pe_empty(
  input [127:0] in_from_east,
  input [127:0] in_from_west,
  input [127:0] in_from_north,
  input [127:0] in_from_south,

  output [127:0] out_to_east,
  output [127:0] out_to_west,
  output [127:0] out_to_north,
  output [127:0] out_to_south,

  input clk,
  input reset
  );


endmodule
